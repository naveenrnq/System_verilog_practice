/*

Encapsulation: Bundles data and methods while restricting direct access to some components, promoting data integrity.

Abstraction: Simplifies complex systems by focusing on essential characteristics and hiding unnecessary details.

Inheritance: Allows classes to inherit attributes and methods from other classes, promoting code reuse and establishing relationships.

Polymorphism: Enables methods to behave differently based on the object type, allowing a unified interface for different implementations.

*/

